module h_rom_l(addr,dout,RisingTone);
input[5:0] addr;
input RisingTone;
output reg[15:0] dout;

always @(*)
begin
   if(~RisingTone)
	   case(addr)
		6'b111111: dout = 16'b1111111111010111;
		6'b111110: dout = 16'b1111111110011000;
		6'b111101: dout = 16'b1111111110001100;
		6'b111100: dout = 16'b1111111111001000;
		6'b111011: dout = 16'b0000000001000011;
		6'b111010: dout = 16'b0000000011000110;
		6'b111001: dout = 16'b0000000011110010;
		6'b111000: dout = 16'b0000000001111010;
		6'b110111: dout = 16'b1111111101101011;
		6'b110110: dout = 16'b1111111001001110;
		6'b110101: dout = 16'b1111110111110111;
		6'b110100: dout = 16'b1111111011111111;
		6'b110011: dout = 16'b0000000100110001;
		6'b110010: dout = 16'b0000001101100010;
		6'b110001: dout = 16'b0000001111110101;
		6'b110000: dout = 16'b0000000111101001;
		6'b101111: dout = 16'b1111110111001000;
		6'b101110: dout = 16'b1111100111001100;
		6'b101101: dout = 16'b1111100011010110;
		6'b101100: dout = 16'b1111110010010011;
		6'b101011: dout = 16'b0000001111110100;
		6'b101010: dout = 16'b0000101100001011;
		6'b101001: dout = 16'b0000110011010001;
		6'b101000: dout = 16'b0000011000110010;
		6'b100111: dout = 16'b1111100010110101;
		6'b100110: dout = 16'b1110101011111111;
		6'b100101: dout = 16'b1110011001111001;
		6'b100100: dout = 16'b1111001011000110;
		6'b100011: dout = 16'b0001000101010011;
		6'b100010: dout = 16'b0011101101011111;
		6'b100001: dout = 16'b0110001111011101;
		6'b100000: dout = 16'b0111110010101010;
		6'b011111: dout = 16'b0111110010101010;
		6'b011110: dout = 16'b0110001111011101;
		6'b011101: dout = 16'b0011101101011111;
		6'b011100: dout = 16'b0001000101010011;
		6'b011011: dout = 16'b1111001011000110;
		6'b011010: dout = 16'b1110011001111001;
		6'b011001: dout = 16'b1110101011111111;
		6'b011000: dout = 16'b1111100010110101;
		6'b010111: dout = 16'b0000011000110010;
		6'b010110: dout = 16'b0000110011010001;
		6'b010101: dout = 16'b0000101100001011;
		6'b010100: dout = 16'b0000001111110100;
		6'b010011: dout = 16'b1111110010010011;
		6'b010010: dout = 16'b1111100011010110;
		6'b010001: dout = 16'b1111100111001100;
		6'b010000: dout = 16'b1111110111001000;
		6'b001111: dout = 16'b0000000111101001;
		6'b001110: dout = 16'b0000001111110101;
		6'b001101: dout = 16'b0000001101100010;
		6'b001100: dout = 16'b0000000100110001;
		6'b001011: dout = 16'b1111111011111111;
		6'b001010: dout = 16'b1111110111110111;
		6'b001001: dout = 16'b1111111001001110;
		6'b001000: dout = 16'b1111111101101011;
		6'b000111: dout = 16'b0000000001111010;
		6'b000110: dout = 16'b0000000011110010;
		6'b000101: dout = 16'b0000000011000110;
		6'b000100: dout = 16'b0000000001000011;
		6'b000011: dout = 16'b1111111111001000;
		6'b000010: dout = 16'b1111111110001100;
		6'b000001: dout = 16'b1111111110011000;
		6'b000000: dout = 16'b1111111111010111;
	   endcase
	else
	   case(addr)
		6'b111111: dout = 16'b1111111111100010;
		6'b111110: dout = 16'b1111111110110010;
		6'b111101: dout = 16'b1111111110101001;
		6'b111100: dout = 16'b1111111111010110;
		6'b111011: dout = 16'b0000000000110011;
		6'b111010: dout = 16'b0000000010010100;
		6'b111001: dout = 16'b0000000010110101;
		6'b111000: dout = 16'b0000000001011100;
		6'b110111: dout = 16'b1111111110010001;
		6'b110110: dout = 16'b1111111010111011;
		6'b110101: dout = 16'b1111111001111001;
		6'b110100: dout = 16'b1111111100111111;
		6'b110011: dout = 16'b0000000011100100;
		6'b110010: dout = 16'b0000001010001001;
		6'b110001: dout = 16'b0000001011111000;
		6'b110000: dout = 16'b0000000101101111;
		6'b101111: dout = 16'b1111111001010110;
		6'b101110: dout = 16'b1111101101011001;
		6'b101101: dout = 16'b1111101010100000;
		6'b101100: dout = 16'b1111110101101110;
		6'b101011: dout = 16'b0000001011110111;
		6'b101010: dout = 16'b0000100001001000;
		6'b101001: dout = 16'b0000100110011100;
		6'b101000: dout = 16'b0000010010100110;
		6'b100111: dout = 16'b1111101010000111;
		6'b100110: dout = 16'b1111000000111111;
		6'b100101: dout = 16'b1110110011011010;
		6'b100100: dout = 16'b1111011000010100;
		6'b100011: dout = 16'b0000110011111110;
		6'b100010: dout = 16'b0010110010000111;
		6'b100001: dout = 16'b0100101011100110;
		6'b100000: dout = 16'b0101110110000000;
		6'b011111: dout = 16'b0101110110000000;
		6'b011110: dout = 16'b0100101011100110;
		6'b011101: dout = 16'b0010110010000111;
		6'b011100: dout = 16'b0000110011111110;
		6'b011011: dout = 16'b1111011000010100;
		6'b011010: dout = 16'b1110110011011010;
		6'b011001: dout = 16'b1111000000111111;
		6'b011000: dout = 16'b1111101010000111;
		6'b010111: dout = 16'b0000010010100110;
		6'b010110: dout = 16'b0000100110011100;
		6'b010101: dout = 16'b0000100001001000;
		6'b010100: dout = 16'b0000001011110111;
		6'b010011: dout = 16'b1111110101101110;
		6'b010010: dout = 16'b1111101010100000;
		6'b010001: dout = 16'b1111101101011001;
		6'b010000: dout = 16'b1111111001010110;
		6'b001111: dout = 16'b0000000101101111;
		6'b001110: dout = 16'b0000001011111000;
		6'b001101: dout = 16'b0000001010001001;
		6'b001100: dout = 16'b0000000011100100;
		6'b001011: dout = 16'b1111111100111111;
		6'b001010: dout = 16'b1111111001111001;
		6'b001001: dout = 16'b1111111010111011;
		6'b001000: dout = 16'b1111111110010001;
		6'b000111: dout = 16'b0000000001011100;
		6'b000110: dout = 16'b0000000010110101;
		6'b000101: dout = 16'b0000000010010100;
		6'b000100: dout = 16'b0000000000110011;
		6'b000011: dout = 16'b1111111111010110;
		6'b000010: dout = 16'b1111111110101001;
		6'b000001: dout = 16'b1111111110110010;
		6'b000000: dout = 16'b1111111111100010;
	   endcase
end

endmodule