module h_rom_h(addr,dout,mode);
input mode;
input[4:0] addr;
output reg[15:0] dout;

always @(*)begin

		if(mode) begin
		case(addr)
			5'b00000: dout = 16'b1111111111011111;
5'b00001: dout = 16'b1111111111001101;
5'b00010: dout = 16'b1111111110101100;
5'b00011: dout = 16'b1111111101111010;
5'b00100: dout = 16'b1111111100110111;
5'b00101: dout = 16'b1111111011110000;
5'b00110: dout = 16'b1111111010110101;
5'b00111: dout = 16'b1111111010100001;
5'b01000: dout = 16'b1111111011010100;
5'b01001: dout = 16'b1111111101110111;
5'b01010: dout = 16'b0000000010111000;
5'b01011: dout = 16'b0000001011011001;
5'b01100: dout = 16'b0000011001001101;
5'b01101: dout = 16'b0000110000101111;
5'b01110: dout = 16'b0001100010010001;
5'b01111: dout = 16'b0101000010011001;
5'b10000: dout = 16'b1010111101100111;
5'b10001: dout = 16'b1110011101101111;
5'b10010: dout = 16'b1111001111010001;
5'b10011: dout = 16'b1111100110110011;
5'b10100: dout = 16'b1111110100100111;
5'b10101: dout = 16'b1111111101001000;
5'b10110: dout = 16'b0000000010001001;
5'b10111: dout = 16'b0000000100101100;
5'b11000: dout = 16'b0000000101011111;
5'b11001: dout = 16'b0000000101001011;
5'b11010: dout = 16'b0000000100010000;
5'b11011: dout = 16'b0000000011001001;
5'b11100: dout = 16'b0000000010000110;
5'b11101: dout = 16'b0000000001010100;
5'b11110: dout = 16'b0000000000110011;
5'b11111: dout = 16'b0000000000100001;
endcase

		end
		else begin
		case(addr)
/*400hz
			5'b00000: dout = 16'b0000000000100101;
5'b00001: dout = 16'b0000000000101111;
5'b00010: dout = 16'b0000000001000101;
5'b00011: dout = 16'b0000000001101100;
5'b00100: dout = 16'b0000000010100111;
5'b00101: dout = 16'b0000000011111011;
5'b00110: dout = 16'b0000000101101111;
5'b00111: dout = 16'b0000001000001001;
5'b01000: dout = 16'b0000001011010100;
5'b01001: dout = 16'b0000001111011111;
5'b01010: dout = 16'b0000010101000110;
5'b01011: dout = 16'b0000011100111100;
5'b01100: dout = 16'b0000101000101101;
5'b01101: dout = 16'b0000111100111001;
5'b01110: dout = 16'b0001101010000010;
5'b01111: dout = 16'b0101000101000100;
5'b10000: dout = 16'b1010111010111100;
5'b10001: dout = 16'b1110010101111110;
5'b10010: dout = 16'b1111000011000111;
5'b10011: dout = 16'b1111010111010011;
5'b10100: dout = 16'b1111100011000100;
5'b10101: dout = 16'b1111101010111010;
5'b10110: dout = 16'b1111110000100001;
5'b10111: dout = 16'b1111110100101100;
5'b11000: dout = 16'b1111110111110111;
5'b11001: dout = 16'b1111111010010001;
5'b11010: dout = 16'b1111111100000101;
5'b11011: dout = 16'b1111111101011001;
5'b11100: dout = 16'b1111111110010100;
5'b11101: dout = 16'b1111111110111011;
5'b11110: dout = 16'b1111111111010001;
5'b11111: dout = 16'b1111111111011011;*/

			

			//200hz
			5'b00000: dout = 16'b0000000000110001;
5'b00001: dout = 16'b0000000000111100;
5'b00010: dout = 16'b0000000001010101;
5'b00011: dout = 16'b0000000010000000;
5'b00100: dout = 16'b0000000011000001;
5'b00101: dout = 16'b0000000100011100;
5'b00110: dout = 16'b0000000110010101;
5'b00111: dout = 16'b0000001000110011;
5'b01000: dout = 16'b0000001100000000;
5'b01001: dout = 16'b0000010000001100;
5'b01010: dout = 16'b0000010101110010;
5'b01011: dout = 16'b0000011101100011;
5'b01100: dout = 16'b0000101001001110;
5'b01101: dout = 16'b0000111101010011;
5'b01110: dout = 16'b0001101010010010;
5'b01111: dout = 16'b0101000101001010;
5'b10000: dout = 16'b1010111010110110;
5'b10001: dout = 16'b1110010101101110;
5'b10010: dout = 16'b1111000010101101;
5'b10011: dout = 16'b1111010110110010;
5'b10100: dout = 16'b1111100010011101;
5'b10101: dout = 16'b1111101010001110;
5'b10110: dout = 16'b1111101111110100;
5'b10111: dout = 16'b1111110100000000;
5'b11000: dout = 16'b1111110111001101;
5'b11001: dout = 16'b1111111001101011;
5'b11010: dout = 16'b1111111011100100;
5'b11011: dout = 16'b1111111100111111;
5'b11100: dout = 16'b1111111110000000;
5'b11101: dout = 16'b1111111110101011;
5'b11110: dout = 16'b1111111111000100;
5'b11111: dout = 16'b1111111111001111;

		/*	0 : dout=16'd65515;
			1 : dout=16'd65512;
			2 : dout=16'd65504;
			3 : dout=16'd65491;
			4 : dout=16'd65474;
			5 : dout=16'd65452;
			6 : dout=16'd65428;
			7 : dout=16'd65403;
			8 : dout=16'd65376;
			9 : dout=16'd65351;
			10: dout=16'd65326;
			11: dout=16'd65305;
			12: dout=16'd65287;
			13: dout=16'd65274;
			14: dout=16'd65266;
			15: dout=16'd32474;*/

			

			/*5'b00000: dout = 16'b1111111111110010;
			5'b00001: dout = 16'b0000000000010001;
			5'b00010: dout = 16'b0000000001000000;
			5'b00011: dout = 16'b0000000010000011;
			5'b00100: dout = 16'b0000000011000011;
			5'b00101: dout = 16'b0000000011010000;
			5'b00110: dout = 16'b0000000001101100;
			5'b00111: dout = 16'b1111111101101011;
			5'b01000: dout = 16'b1111110111010110;
			5'b01001: dout = 16'b1111110000001000;
			5'b01010: dout = 16'b1111101010110000;
			5'b01011: dout = 16'b1111101010111101;
			5'b01100: dout = 16'b1111110101010010;
			5'b01101: dout = 16'b0000001111111001;
			5'b01110: dout = 16'b0001001011001101;
			5'b01111: dout = 16'b0100111010000110;
			5'b10000: dout = 16'b1011000101111010;
			5'b10001: dout = 16'b1110110100110011;
			5'b10010: dout = 16'b1111110000000111;
			5'b10011: dout = 16'b0000001010101110;
			5'b10100: dout = 16'b0000010101000011;
			5'b10101: dout = 16'b0000010101010000;
			5'b10110: dout = 16'b0000001111111000;
			5'b10111: dout = 16'b0000001000101010;
			5'b11000: dout = 16'b0000000010010101;
			5'b11001: dout = 16'b1111111110010100;
			5'b11010: dout = 16'b1111111100110000;
			5'b11011: dout = 16'b1111111100111101;
			5'b11100: dout = 16'b1111111101111101;
			5'b11101: dout = 16'b1111111111000000;
			5'b11110: dout = 16'b1111111111101111;
			5'b11111: dout = 16'b0000000000001110;*/
				/*5'b00000: dout = 16'b1111111111011111;
				5'b00001: dout = 16'b1111111111001101;
				5'b00010: dout = 16'b1111111110101100;
				5'b00011: dout = 16'b1111111101111010;
				5'b00100: dout = 16'b1111111100110111;
				5'b00101: dout = 16'b1111111011110000;
				5'b00110: dout = 16'b1111111010110101;
				5'b00111: dout = 16'b1111111010100001;
				5'b01000: dout = 16'b1111111011010100;
				5'b01001: dout = 16'b1111111101110111;
				5'b01010: dout = 16'b0000000010111000;
				5'b01011: dout = 16'b0000001011011001;
				5'b01100: dout = 16'b0000011001001101;
				5'b01101: dout = 16'b0000110000101111;
				5'b01110: dout = 16'b0001100010010001;
				5'b01111: dout = 16'b0101000010011001;
				5'b10000: dout = 16'b1010111101100111;
				5'b10001: dout = 16'b1110011101101111;
				5'b10010: dout = 16'b1111001111010001;
				5'b10011: dout = 16'b1111100110110011;
				5'b10100: dout = 16'b1111110100100111;
				5'b10101: dout = 16'b1111111101001000;
				5'b10110: dout = 16'b0000000010001001;
				5'b10111: dout = 16'b0000000100101100;
				5'b11000: dout = 16'b0000000101011111;
				5'b11001: dout = 16'b0000000101001011;
				5'b11010: dout = 16'b0000000100010000;
				5'b11011: dout = 16'b0000000011001001;
				5'b11100: dout = 16'b0000000010000110;
				5'b11101: dout = 16'b0000000001010100;
				5'b11110: dout = 16'b0000000000110011;
				5'b11111: dout = 16'b0000000000100001;*/
			endcase
			
		end
			
end

endmodule